module codemem ();

endmodule