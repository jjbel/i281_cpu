module User_Code_Low(b0I,b1I,b2I,b3I,b4I,b5I,b6I,b7I,b8I,b9I,b10I,b11I,b12I,b13I,b14I,b15I);

output [16:0] b0I;
output [16:0] b1I;
output [16:0] b2I;
output [16:0] b3I;
output [16:0] b4I;
output [16:0] b5I;
output [16:0] b6I;
output [16:0] b7I;
output [16:0] b8I;
output [16:0] b9I;
output [16:0] b10I;
output [16:0] b11I;
output [16:0] b12I;
output [16:0] b13I;
output [16:0] b14I;
output [16:0] b15I;

assign b0I[16:0] = 17'b0_0011_00_00_00000000;
assign b1I[16:0] = 17'b0_1000_11_00_00001000;
assign b2I[16:0] = 17'b0_0011_01_00_00000000;
assign b3I[16:0] = 17'b0_1101_00_11_00000000;
assign b4I[16:0] = 17'b0_1111_00_11_00001110;
assign b5I[16:0] = 17'b0_1000_11_00_00001000;
assign b6I[16:0] = 17'b0_0110_11_00_00000000;
assign b7I[16:0] = 17'b0_1101_01_11_00000000;
assign b8I[16:0] = 17'b0_1111_00_11_00001000;
assign b9I[16:0] = 17'b0_1001_10_01_00000000;
assign b10I[16:0] = 17'b0_1001_11_01_00000001;
assign b11I[16:0] = 17'b0_1101_11_10_00000000;
assign b12I[16:0] = 17'b0_1111_00_11_00000010;
assign b13I[16:0] = 17'b0_1011_11_01_00000000;
assign b14I[16:0] = 17'b0_1011_10_01_00000001;
assign b15I[16:0] = 17'b0_0101_01_00_00000001;
endmodule
