/*
i281 Top Level Entity
*/

//module includes
`include "ALU/alu.v"
`include "Code Memory/codemem.v"
`include "Control Logic/controllogic.v"
`include "Data Memory/datamem.v"
`include "Flags/flags.v"
`include "OpCode Decoder/opcodedec.v"
`include "PC/pc.v"
`include "Registers/register.v"

//