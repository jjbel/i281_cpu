module BIOS_Hardcoded_High(b0I,b1I,b2I,b3I,b4I,b5I,b6I,b7I,b8I,b9I,b10I,b11I,b12I,b13I,b14I,b15I);
//BIOS v17.0 1/3/2019
//author: Alexander Stoytchev
output [16:0] b0I;
output [16:0] b1I;
output [16:0] b2I;
output [16:0] b3I;
output [16:0] b4I;
output [16:0] b5I;
output [16:0] b6I;
output [16:0] b7I;
output [16:0] b8I;
output [16:0] b9I;
output [16:0] b10I;
output [16:0] b11I;
output [16:0] b12I;
output [16:0] b13I;
output [16:0] b14I;
output [16:0] b15I;

//multicycle flag added as MSB

assign b0I[16:0] = 17'b0_0000_00_00_00000000;
assign b1I[16:0] = 17'b0_0000_00_00_00000000;
assign b2I[16:0] = 17'b0_0000_00_00_00000000;
assign b3I[16:0] = 17'b0_0000_00_00_00000000;
assign b4I[16:0] = 17'b0_0000_00_00_00000000;
assign b5I[16:0] = 17'b0_0000_00_00_00000000;
assign b6I[16:0] = 17'b0_0000_00_00_00000000;
assign b7I[16:0] = 17'b0_0000_00_00_00000000;
assign b8I[16:0] = 17'b0_0000_00_00_00000000;
assign b9I[16:0] = 17'b0_0000_00_00_00000000;
assign b10I[16:0] = 17'b0_0000_00_00_00000000;
assign b11I[16:0] = 17'b0_0000_00_00_00000000;
assign b12I[16:0] = 17'b0_0000_00_00_00000000;
assign b13I[16:0] = 17'b0_0000_00_00_00000000;
assign b14I[16:0] = 17'b0_0000_00_00_00000000;
assign b15I[16:0] = 17'b0_0000_00_00_00000000;

endmodule